module testeINOUT(entrada);

    inout entrada;

endmodule